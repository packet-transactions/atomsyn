module counter(
    //--------------------------------------------------------------------------
    // Global signals
    //--------------------------------------------------------------------------
    clk,

    //--------------------------------------------------------------------------
    // Input interface
    //--------------------------------------------------------------------------
    i__inc,

    //--------------------------------------------------------------------------
    // Output interface
    //--------------------------------------------------------------------------
    o__count__next
);

//------------------------------------------------------------------------------
// Parameters
//------------------------------------------------------------------------------
parameter COUNT_WIDTH                   = 3;
parameter INIT_VALUE                    = 1'b0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Global signals
//------------------------------------------------------------------------------
input  logic                            clk;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Input interface
//------------------------------------------------------------------------------
input  logic                            i__inc;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output interface
//------------------------------------------------------------------------------
output logic [COUNT_WIDTH-1:0]          o__count__next;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Internal signals
//------------------------------------------------------------------------------
logic [COUNT_WIDTH-1:0]                 r__count__pff;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Count logic
//------------------------------------------------------------------------------
always_comb
begin
    o__count__next = r__count__pff;

    if(i__inc == 1'b1)
    begin
        if(r__count__pff == 7)
        begin
            o__count__next = '0;
        end
        else
        begin
            o__count__next = r__count__pff + 1'b1;
        end
    end
end

always_ff @ (posedge clk)
begin
    r__count__pff <= o__count__next;
end
//------------------------------------------------------------------------------

endmodule
